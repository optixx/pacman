-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity PACROM_5E is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(11 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of PACROM_5E is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S4
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (3 downto 0);
      ADDR  : in  std_logic_vector (11 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (3 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(11 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(11 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "00445764023999F602644573037FDD91000277000011FF11013446310CE311EC";
    attribute INIT_01 of inst : label is "066445760007F800013644400EF999F607755550023111FE001367700CC44FF4";
    attribute INIT_02 of inst : label is "077444730FF999F6013646310FF444FF0374447300999BEC037544300699DD76";
    attribute INIT_03 of inst : label is "077444440FF888800077444400FF9991077446310FF113EC013644620CE31132";
    attribute INIT_04 of inst : label is "00133100008CC80000133100008CC80000011000000880000001100000088000";
    attribute INIT_05 of inst : label is "0000000000000000000000000000000037FFFF73CEFFFFEC37FFFF73CEFFFFEC";
    attribute INIT_06 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_07 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_08 of inst : label is "0002377F00000888FFFEC000880000000000133300088CCE33100000EFFF7000";
    attribute INIT_09 of inst : label is "00DE0DE00000000000DE0DE00000000000000000066000000000000000000000";
    attribute INIT_0A of inst : label is "FFCCF700FF00FF00F700FFCCFF00FF00001DDDDD00FFBBBBFFCCCCF7FF0000FF";
    attribute INIT_0B of inst : label is "0000000000000000F7000000FE000000007FCCCC00EF33337FCCCCCCEF333333";
    attribute INIT_0C of inst : label is "0089BFD8046222EC04C99BF606EEAA220004FF000022EE2203788C7308C622C8";
    attribute INIT_0D of inst : label is "0CC89BEC000EE000037D99900CE222EC0EEAAAB1046222EC0136CFF008888EE8";
    attribute INIT_0E of inst : label is "0001110000000000000012480248000006F999F7002226C806FB99600C22AAEC";
    attribute INIT_0F of inst : label is "F0000000F1111111F8888888F00000000000000F1111111F8888888F0000000F";
    attribute INIT_10 of inst : label is "037C88C408C622640FF999F60EE222EC037C8C730EE888EE0000000000000000";
    attribute INIT_11 of inst : label is "037C899908C622EE0FF999980EE0000000FF999800EE22220FF88C730EE226C8";
    attribute INIT_12 of inst : label is "0FF136C80EE8CE62000000FF046222EC0088FF880022EE220FF111FF0EE000EE";
    attribute INIT_13 of inst : label is "07F888F70CE222EC0FF731FF0EE08CEE0FF737FF0EE080EE00FF000000EE2222";
    attribute INIT_14 of inst : label is "06F99D50046222EC0FF889F70EE8CE6207F888F70CE2AECA0FF888F70EE88880";
    attribute INIT_15 of inst : label is "0FF131FF0EEC8CEE0FF101FF008CEC800FF000FF0CE222EC0088FF880000EE00";
    attribute INIT_16 of inst : label is "0003FEC0002800000889BFEC06EEA22200EF11FE0000EE000CE737EC06EC8CE6";
    attribute INIT_17 of inst : label is "200000004000000032201222E0002AAA32221022E8880000349AA843C295512C";
    attribute INIT_18 of inst : label is "0EEEEEEE00000000033330000FFFFF730000000E000000000000000000000001";
    attribute INIT_19 of inst : label is "00000EEE000000000000033300000FFFEEEEEEEE0000000033100000FFFF7733";
    attribute INIT_1A of inst : label is "000EEEEE0000000000033331000FFFFFEEEEEEEE0000000000000000F7733333";
    attribute INIT_1B of inst : label is "000000000000000000000000000000000226EEEE000000000000000000000013";
    attribute INIT_1C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "EAAA90784222C0C288AD80784222C0C2004F0078002E20C20000000000000000";
    attribute INIT_21 of inst : label is "00000068000000264F0078872E20C22C870788702C0C22C0C88BC07800E000C2";
    attribute INIT_22 of inst : label is "000000EA00000042AD80788722C0C22C000000880000004289607887A220C22C";
    attribute INIT_23 of inst : label is "0000000000000000870000002C000000078870780C22C0C2AA90788722C0C22C";
    attribute INIT_24 of inst : label is "00EFFF8700000008F3FF7000CCCC800000000000001332110000000000000000";
    attribute INIT_25 of inst : label is "008EFFFF0000088CFFEE80008800000000000003007FF7730000000077FF7000";
    attribute INIT_26 of inst : label is "00EFFFFF00088CCCFFFFFE00CCC88000000000010013777F0000000077773100";
    attribute INIT_27 of inst : label is "003FC7FF00C88888FFFFF300EE888C00000001120001FCBF21100000FFFF1000";
    attribute INIT_28 of inst : label is "00CFFFFF00008CC8FFFFFC00CCC800000001110000FFFFF701110000FFFFF700";
    attribute INIT_29 of inst : label is "0000EA15000000485B1C400002480000000004220000023232200000C1120000";
    attribute INIT_2A of inst : label is "008CEF8F0000000C8FEC8000000000000000000000F31130000000003113F000";
    attribute INIT_2B of inst : label is "000000F0000000C2D8000000C800000000000000000000100000000010000000";
    attribute INIT_2C of inst : label is "FFFF9930FFFFFFF003FFFF990FFFFFFF00000000FF77310000000000001377FF";
    attribute INIT_2D of inst : label is "000000000000000000000000000000000CC808C0000000000C808CC000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "F00F0000F00F00000000F00F0000F00F03448999F0078000999844300008700F";
    attribute INIT_35 of inst : label is "F00E1000F00008880001E00F8880000FF00E10000C2219990001E00F999122C0";
    attribute INIT_36 of inst : label is "99999999000000009999999900000000F0000111F00780001110000F0008700F";
    attribute INIT_37 of inst : label is "0000000088888888000000008888888800000000999999990000000099999999";
    attribute INIT_38 of inst : label is "000000000344888800000000888844300C22111100000000111122C000000000";
    attribute INIT_39 of inst : label is "0000000000003488000000008843000011111111000000001111111100000000";
    attribute INIT_3A of inst : label is "0000C21100000000112C0000000000000000F0000000F000000F0000000F0000";
    attribute INIT_3B of inst : label is "0000F11900000000911F000000000000000000000000F88900000000988F0000";
    attribute INIT_3C of inst : label is "11100000000870000000011100078000000000009999999F00000000F9999999";
    attribute INIT_3D of inst : label is "000000000000348800000000884300000001E00088800000000E100000000888";
    attribute INIT_3E of inst : label is "999888880008700088888999000780000000C21100000000112C000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S4
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0000",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "00445764023999F602644573037FDD91000277000011FF11013446310CE311EC";
    attribute INIT_01 of inst : label is "066445760007F800013644400EF999F607755550023111FE001367700CC44FF4";
    attribute INIT_02 of inst : label is "077444730FF999F6013646310FF444FF0374447300999BEC037544300699DD76";
    attribute INIT_03 of inst : label is "077444440FF888800077444400FF9991077446310FF113EC013644620CE31132";
    attribute INIT_04 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_05 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_06 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_07 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_08 of inst : label is "0002377F00000888FFFEC000880000000000133300088CCE33100000EFFF7000";
    attribute INIT_09 of inst : label is "00DE0DE00000000000DE0DE00000000000000000066000000000000000000000";
    attribute INIT_0A of inst : label is "FFCCF700FF00FF00F700FFCCFF00FF00001DDDDD00FFBBBBFFCCCCF7FF0000FF";
    attribute INIT_0B of inst : label is "0000000000000000F7000000FE000000007FCCCC00EF33337FCCCCCCEF333333";
    attribute INIT_0C of inst : label is "0089BFD8046222EC04C99BF606EEAA220004FF000022EE2203788C7308C622C8";
    attribute INIT_0D of inst : label is "0CC89BEC000EE000037D99900CE222EC0EEAAAB1046222EC0136CFF008888EE8";
    attribute INIT_0E of inst : label is "0001110000000000000012480248000006F999F7002226C806FB99600C22AAEC";
    attribute INIT_0F of inst : label is "F0000000F1111111F8888888F00000000000000F1111111F8888888F0000000F";
    attribute INIT_10 of inst : label is "037C88C408C622640FF999F60EE222EC037C8C730EE888EE0000000000000000";
    attribute INIT_11 of inst : label is "037C899908C622EE0FF999980EE0000000FF999800EE22220FF88C730EE226C8";
    attribute INIT_12 of inst : label is "0FF136C80EE8CE62000000FF046222EC0088FF880022EE220FF111FF0EE000EE";
    attribute INIT_13 of inst : label is "07F888F70CE222EC0FF731FF0EE08CEE0FF737FF0EE080EE00FF000000EE2222";
    attribute INIT_14 of inst : label is "06F99D50046222EC0FF889F70EE8CE6207F888F70CE2AECA0FF888F70EE88880";
    attribute INIT_15 of inst : label is "0FF131FF0EEC8CEE0FF101FF008CEC800FF000FF0CE222EC0088FF880000EE00";
    attribute INIT_16 of inst : label is "0003FEC0002800000889BFEC06EEA22200EF11FE0000EE000CE737EC06EC8CE6";
    attribute INIT_17 of inst : label is "200000004000000032201222E0002AAA32221022E8880000349AA843C295512C";
    attribute INIT_18 of inst : label is "0EEEEEEE00000000033330000FFFFF7300000000000000000000000000000000";
    attribute INIT_19 of inst : label is "00000EEE000000000000033300000FFFEEEEEEEE0000000033100000FFFF7733";
    attribute INIT_1A of inst : label is "000EEEEE0000000000033331000FFFFFEEEEEEEE0000000000000000F7733333";
    attribute INIT_1B of inst : label is "000000000000000000000000000000000226EEEC000000000000000000000013";
    attribute INIT_1C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "EAAA90784222C0C288AD80784222C0C2004F0078002E20C20000000000000000";
    attribute INIT_21 of inst : label is "00000068000000264F0078872E20C22C870788702C0C22C0C88BC07800E000C2";
    attribute INIT_22 of inst : label is "000000EA00000042AD80788722C0C22C000000880000004289607887A220C22C";
    attribute INIT_23 of inst : label is "0000000000000000870000002C000000078870780C22C0C2AA90788722C0C22C";
    attribute INIT_24 of inst : label is "00042000000000001C00000008000000000000000000012400113300892C0000";
    attribute INIT_25 of inst : label is "00004014000000000180000000000000000011130002098D111000008A040000";
    attribute INIT_26 of inst : label is "00000000000000000000000000000000000000010000004E1331100048880000";
    attribute INIT_27 of inst : label is "0000000000066666000000006666600000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000002C00000000000000000001000000082000000000000000";
    attribute INIT_29 of inst : label is "000EB5EF00008C86A5E7BE00EC848000000000000000356D00000000BF653000";
    attribute INIT_2A of inst : label is "00008C8F0000000C8C8000000000000000000001000337FF00000000F7330000";
    attribute INIT_2B of inst : label is "000000F0000000C2D8000000C8000000000011220000EEFE21100000FEE00000";
    attribute INIT_2C of inst : label is "FF106730FFFFFFF003FF10670FFFFFFF00000000FF76210000000000001376EF";
    attribute INIT_2D of inst : label is "000000000000000000000000000000000CC808C0000000000C808CC000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000066666666000000006666666600000000000000000000000000000000";
    attribute INIT_34 of inst : label is "FFFF0000FFFF00000000FFFF0000FFFF0377FFFFFFFF8000FFFF77300008FFFF";
    attribute INIT_35 of inst : label is "FFFF1000FFFFFFFF0001FFFFFFFFFFFFFFFF10000CEEFFFF0001FFFFFFFFEEC0";
    attribute INIT_36 of inst : label is "FFFFFFFF00000000FFFFFFFF00000000FFFFFFFFFFFF8000FFFFFFFF0008FFFF";
    attribute INIT_37 of inst : label is "00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF";
    attribute INIT_38 of inst : label is "000000000377FFFF00000000FFFF77300CEEFFFF00000000FFFFEEC000000000";
    attribute INIT_39 of inst : label is "00000000000037FF00000000FF730000FFFFFFFF00000000FFFFFFFF00000000";
    attribute INIT_3A of inst : label is "0000CEFF00000000FFEC0000000000000000FFFF0000FFFFFFFF0000FFFF0000";
    attribute INIT_3B of inst : label is "0000FFFF00000000FFFF000000000000000000000000FFFF00000000FFFF0000";
    attribute INIT_3C of inst : label is "FFFFFFFF0008FFFFFFFFFFFFFFFF800000000000FFFFFFFF00000000FFFFFFFF";
    attribute INIT_3D of inst : label is "00000000000037FF00000000FF7300000001FFFFFFFFFFFFFFFF1000FFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFF0008FFFFFFFFFFFFFFFF80000000CEFF00000000FFEC000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S4
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0000",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
